package CONSTANTS is
   constant NB : integer := 11; -- Number of bits
   constant NT : integer := 11; -- Number of taps
   constant L : integer := 3; -- Unfolding degree
end CONSTANTS;

